library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use work.common_pack.all;

entity patRecog is
end patRecog
